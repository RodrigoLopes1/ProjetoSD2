--Agora com o fluxo de dados feito, seria necessário só testar numa testbench de verdade, esse é o objetivo dessa entrega
--A testbench tem que gerar os sinais de Rd, Rn, e Rm e outras coisas ai...
