--Vai sair parte 2 tenham fé
