--Vai sair, tenham fé
